* C:\Users\Fariha Rahman\Desktop\PSpice\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Fri Nov 20 14:50:27 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
